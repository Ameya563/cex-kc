module arbiter4( r1, r2, r3, r4, g1, g2, g3, g4, res );
input r1;
input r2;
input r3;
input r4;
input g1;
input g2;
input g3;
input g4;
output res;
wire v1;
wire v2;
wire v3;
wire v4;
wire v5;
wire single;
wire w1;
wire w2;
wire w3;
wire w4;
wire causal;
wire off;
wire x;
assign v1 = (g1 & ~g2 & ~g3 & ~g4);
assign v2 = (g2 & ~g3 & ~g1 & ~g4);
assign v3 = (g3 & ~g1 & ~g2 & ~g4);
assign v4 = (g4 & ~g1 & ~g2 & ~g3);
assign v5 = (~g1 & ~g2 & ~g3 & ~g4);
assign single = (v1 | v2 | v3 | v4 | v5);
assign w1 = (r1 | ~g1);
assign w2 = (r2 | ~g2);
assign w3 = (r3 | ~g3);
assign w4 = (r4 | ~g4);
assign causal = (w1 & w2 & w3 & w4);
assign off = (~r1 & ~r2 & ~r3 & ~r4);
assign x = (~v5 | off);
assign res = (single & causal & x);

endmodule